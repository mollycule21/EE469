module test (input logic x, output logic );'

	assign y = x;
	
endmodule 
