module data_memory();



endmodule
