// 32 regs in RV32i

module reg_file();


endmodule
