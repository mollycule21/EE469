// control signals for alu is defined here

localparam [2:0]ALU_ADD = 3'b000;
localparam [2:0]ALU_SUB = 3'b001;
localparam [2:0]ALU_AND = 3'b010;
localparam [2:0]ALU_OR  = 3'b011;
localparam [2:0]ALU_XOR = 3'b100;
localparam [2:0]ALU_SL  = 3'b101;
localparam [2:0]ALU_SRL = 3'b110;
localparam [2:0]ALU_SRA = 3'b111;
