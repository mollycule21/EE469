module decoder5_32();




endmodule
