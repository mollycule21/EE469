module control_signals;



endmodule
