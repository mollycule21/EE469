module decoder5_32(in, sel, out);
	input logic [4:0]in;
	input logic 



endmodule
